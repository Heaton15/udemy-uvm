`include "uvm_macros.svh"
import uvm_pkg::*;


module tb;
  initial begin
    run_test("test");
  end
endmodule
